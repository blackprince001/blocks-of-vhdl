-- TIPS
    -- place each entity in a different file
    -- current directory of project is always referenced as work.


-- MODELLING STYLES
    -- dataflow: concurrent statements
    -- structural: components and interconnects
    -- behavioural: sequential states (registers, state machines, decoders)
        -- some behavioural descriptions cannot be synthesized!

    -- STRUCTURAL MODELLING

-- precedence of operators
 -- implied precedence

-- Modelling Routing Structures

-- when else structures construct

-- conditional concurrent signal assignment

-- precedence of operators
 -- implied precedence

-- Modelling Routing Structures

-- when else structures construct
-- relational operators and their precedence

-- selective conditional concurrent signal assignment