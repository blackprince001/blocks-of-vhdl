-- test benching

-- waveform viewing or automated checking for observing signal outputs of components
-- or architectures
