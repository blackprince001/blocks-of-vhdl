-- TIPS
    -- place each entity in a different file
    -- current directory of project is always referenced as work.


-- MODELLING STYLES
    -- dataflow: concurrent statements
    -- structural: components and interconnects
    -- behavioural: sequential states (registers, state machines, decoders)
        -- some behavioural descriptions cannot be synthesized!

    -- STRUCTURAL MODELLING