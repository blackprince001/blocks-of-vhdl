-- what is the use if you are only giving me linting
library ieee;
use ieee.std_logic_1164.all;

entity ent is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig : out std_logic
    );
end ent;

architecture rtl of ent is
    
begin

end architecture;